//========================================================================
// Nor Gate-Level Model
//========================================================================

module NorGL
(
  input  a,
  input  b,
  output y
);

  assign y = !( a | b );

endmodule

